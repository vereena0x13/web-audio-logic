module not1(
    input wire a,
    output wire y
);

    assign y = ~a;

endmodule
