module add1(
    input wire [2:0] a,
    output wire [2:0] y
);

    assign y = a + 3'd1;

endmodule
